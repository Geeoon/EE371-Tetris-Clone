module clear_row_data(init_regs, clk, incr_row, row, final_row);
	input logic init_regs, clk, incr_row;
	
	output logic [4:0] row;
	output logic final_row;
	
	always_ff @(posedge clk) begin
			if(init_regs) begin
				row <= 0;
			end
			if (incr_row) begin
				row <= row + 5'b1;
			end
		end //always_ff
		
		assign final_row = (row == 19);
endmodule